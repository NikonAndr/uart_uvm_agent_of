interface uart_if();
    logic tx;
    logic rst;
endinterface : uart_if